--------------------------------------------------------------------------------
-- Module Name: Follow here with one phrase describing module.
--
-- Created by: Daniel C. Nygren
-- Email: dan.nygren@gmail.com
-- Permanent Email: Dan.Nygren@alumni.clemson.edu
--
-- Copyright 2019 by Daniel C. Nygren
--
--   Permission to use and modify this software for any purpose other than
-- its incorporation into a commercial product is hereby granted without fee.
-- Permission to copy and distribute this software only for non-commercial use
-- is also granted without fee, provided that the above copyright notice and
-- this entire permission notice appear in all copies and any supporting
-- documentation. The author makes no representations about the suitability of
-- this software for any purpose. It is provided "as is" without express or
-- implied warranty.
--
--   Start here a paragraph explaining what the module does and how it works.
-- Include a description of module limitations and algorithms.
--
-- CALLING SEQUENCE  (Example with explanation of call parameters)
--
-- EXAMPLES          (Examples of calls)
--
-- TARGET SYSTEM     (System code targeted for)
--
-- DEVELOPED USING   (System code developed on)
--
-- CALLS             (List of modules this routine calls)
--
-- CALLED BY         (List of modules that call this one)
--
-- INPUTS            (Parameters used but not modified, include global and
--                   static data)
--
-- OUTPUTS           (Parameters modified, include global and static data)
--
-- RETURNS           (Type and meaning of return value, if any)
--
-- ERROR HANDLING    (Describe how errors are handled)
--
-- WARNINGS          (1. Describe anything a maintainer should be aware of)
--                   (2. Describe anything a maintainer should be aware of)
--                   (N. Describe anything a maintainer should be aware of)
--------------------------------------------------------------------------------

-- (Delete this explanation from your code.)
-- The below lines are optionally used to aid maintainers by indicating at
-- which point portions of the code intended or likely to be modified end.

-- ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
-- ^^^^^^^^^^ Place code that may need modification above this point. ^^^^^^^^^^
-- ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
