--------------------------------------------------------------------------------
-- Module Name: Follow here with one phrase describing module.
--
-- Created by: Daniel C. Nygren
-- Email: nygren@msss.com
-- Permanent Email: dan.nygren@gmail.com
--
-- Copyright (c) 2001, 2024, Daniel C. Nygren.
--
-- BSD 0-clause license, "Zero Clause BSD", SPDX: 0BSD
--
-- Permission to use, copy, modify, and/or distribute this software for any
-- purpose with or without fee is hereby granted.
--
-- THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES WITH
-- REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF MERCHANTABILITY
-- AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR ANY SPECIAL, DIRECT,
-- INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES WHATSOEVER RESULTING FROM
-- LOSS OF USE, DATA OR PROFITS, WHETHER IN AN ACTION OF CONTRACT, NEGLIGENCE
-- OR OTHER TORTIOUS ACTION, ARISING OUT OF OR IN CONNECTION WITH THE USE OR
-- PERFORMANCE OF THIS SOFTWARE.
--
--   Start here a paragraph explaining what the module does and how it works.
-- Include a description of module limitations and algorithms.
--
-- CALL SEQUENCE  (Example with explanation of call parameters)
--
-- EXAMPLES       (Examples of calls)
--
-- TARGET SYSTEM  (System code targeted for)
--
-- DEVELOPED ON   (System code developed on)
--
-- CALLS          (List of modules this routine calls)
--
-- CALLED BY      (List of modules that call this one)
--
-- INPUTS         (Parameters used but not modified, include global/static data)
--
-- OUTPUTS        (Parameters modified, include global/static data)
--
-- RETURNS        (Type and meaning of return value, if any)
--
-- ERROR HANDLING (Describe how errors are handled)
--
-- SECURE CODING  (List methods used to prevent exploits against this code)
--
-- WARNINGS       (1. Describe anything a maintainer should be aware of)
--                (2. Describe anything a maintainer should be aware of)
--                (N. Describe anything a maintainer should be aware of)
--------------------------------------------------------------------------------

-- (Delete this explanation from your code.)
-- The below lines are optionally used to aid maintainers by indicating at
-- which point portions of the code intended or likely to be modified end.

-- ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
-- ^^^^^^^^^^ Place code that may need modification above this point. ^^^^^^^^^^
-- ^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
